module led_encoder(in, out1, out2, out3, out4);
    input wire[15:0] in;
    output reg[6:0] out1;
    output reg[6:0] out2;
    output reg[6:0] out3;
    output reg[6:0] out4;

    always@(*) begin
        case(in[3:0])
            4'b0000: out1 = 7'b0111111; // 0
            4'b0001: out1 = 7'b0000110; // 1
            4'b0010: out1 = 7'b1011011; // 2
            4'b0011: out1 = 7'b1001111; // 3
            4'b0100: out1 = 7'b1100110; // 4
            4'b0101: out1 = 7'b1101101; // 5
            4'b0110: out1 = 7'b1111101; // 6
            4'b0111: out1 = 7'b0000111; // 7
            4'b1000: out1 = 7'b1111111; // 8
            4'b1001: out1 = 7'b1101111; // 9
            4'b1010: out1 = 7'b1110111; // A
            4'b1011: out1 = 7'b1111100; // b
            4'b1100: out1 = 7'b0111001; // C
            4'b1101: out1 = 7'b1011110; // d
            4'b1110: out1 = 7'b1111001; // E
            4'b1111: out1 = 7'b1110001; // F
        endcase

        case(in[7:4])
            4'b0000: out2 = 7'b0111111; // 0
            4'b0001: out2 = 7'b0000110; // 1
            4'b0010: out2 = 7'b1011011; // 2
            4'b0011: out2 = 7'b1001111; // 3
            4'b0100: out2 = 7'b1100110; // 4
            4'b0101: out2 = 7'b1101101; // 5
            4'b0110: out2 = 7'b1111101; // 6
            4'b0111: out2 = 7'b0000111; // 7
            4'b1000: out2 = 7'b1111111; // 8
            4'b1001: out2 = 7'b1101111; // 9
            4'b1010: out2 = 7'b1110111; // A
            4'b1011: out2 = 7'b1111100; // b
            4'b1100: out2 = 7'b0111001; // C
            4'b1101: out2 = 7'b1011110; // d
            4'b1110: out2 = 7'b1111001; // E
            4'b1111: out2 = 7'b1110001; // F
        endcase

        case(in[11:8])
            4'b0000: out3 = 7'b0111111; // 0
            4'b0001: out3 = 7'b0000110; // 1
            4'b0010: out3 = 7'b1011011; // 2
            4'b0011: out3 = 7'b1001111; // 3
            4'b0100: out3 = 7'b1100110; // 4
            4'b0101: out3 = 7'b1101101; // 5
            4'b0110: out3 = 7'b1111101; // 6
            4'b0111: out3 = 7'b0000111; // 7
            4'b1000: out3 = 7'b1111111; // 8
            4'b1001: out3 = 7'b1101111; // 9
            4'b1010: out3 = 7'b1110111; // A
            4'b1011: out3 = 7'b1111100; // b
            4'b1100: out3 = 7'b0111001; // C
            4'b1101: out3 = 7'b1011110; // d
            4'b1110: out3 = 7'b1111001; // E
            4'b1111: out3 = 7'b1110001; // F
        endcase

        case(in[15:12])
            4'b0000: out4 = 7'b0111111; // 0
            4'b0001: out4 = 7'b0000110; // 1
            4'b0010: out4 = 7'b1011011; // 2
            4'b0011: out4 = 7'b1001111; // 3
            4'b0100: out4 = 7'b1100110; // 4
            4'b0101: out4 = 7'b1101101; // 5
            4'b0110: out4 = 7'b1111101; // 6
            4'b0111: out4 = 7'b0000111; // 7
            4'b1000: out4 = 7'b1111111; // 8
            4'b1001: out4 = 7'b1101111; // 9
            4'b1010: out4 = 7'b1110111; // A
            4'b1011: out4 = 7'b1111100; // b
            4'b1100: out4 = 7'b0111001; // C
            4'b1101: out4 = 7'b1011110; // d
            4'b1110: out4 = 7'b1111001; // E
            4'b1111: out4 = 7'b1110001; // F
        endcase
    end
endmodule
