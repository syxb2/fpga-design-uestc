module decoder_3_8(a, b, c, out);
    input a,b,c;  //端口定义
    output reg [7:0] out;//对out定义为1个8位的数据
    //always块描述的信号赋值，被赋值对象必须定义为reg
    // reg [7:0] out; //定义out为1个8位的寄存器

    always @(*) begin
        out[0] = !a && !b && !c;
        out[1] = !a && !b && c;
        out[2] = !a && b && !c;
        out[3] = !a && b && c;
        out[4] = a && !b && !c;
        out[5] = a && !b && c;
        out[6] = a && b && !c;
        out[7] = a && b && c;
        //一个等价的写法是always @(a, b, c),其中的*表示通配符
        //always表示一个语法块
        // case ({a,b,c}) //里面的大括号内容：{a,b.c}表示一个3位的信号这种操作叫做拼接
        //     3'b000: out = 8'b0000_0001;  //b表示binary 二进制，3'b000，表示一个3位的二进制信号，值为000
        //     3'b001: out = 8'b00000010;  //还有常用的格式，比如 d是十进制，3'd5，表示一个3位的十进制信号，值为5和3'b101完全等价
        //     3'b010: out = 8'b00000100;  //h是十六进制 
        //     3'b011: out = 8'b00001000;   //o是八进制符号
        //     3'b100: out = 8'b00010000;
        //     3'b101: out = 8'b00100000;
        //     3'b110: out = 8'b01000000;
        //     3'b111: out = 8'b10000000;
        // endcase
    end
    //一个拼接的例子
    //wire [3:0]d;
    //assign d = {a,1'b0,b,c};
    //拼接了一个四位的信号，其中第一位是a，第二位是0，第三位是b，第四位是c
endmodule

