module control_unit (
    input wire z,
    input wire [3:0] op,
    output reg m2reg,
    output reg PCsrc,
    output reg wmem,
    output reg [2:0] aluc,
    output reg alusrc,
    output reg wreg
);
    
endmodule