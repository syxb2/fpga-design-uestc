/**
 * @brief 控制模块
 */
module ctrl(
    input wire clk,
    input wire rst_n,
    input wire rx,
    output reg [7:0] data,
    output reg rxd
);

endmodule
